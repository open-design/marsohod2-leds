module hexLEDDriver(input [7:0] value, output [6:0] out);

    reg [6:0] segments;

    always @(value)
        begin
            case (value)
                8'h0:   segments = 7'h3F;
                8'h1:   segments = 7'h06;
                8'h2:   segments = 7'h5B;
                8'h3:   segments = 7'h4F;
                8'h4:   segments = 7'h66;
                8'h5:   segments = 7'h6D;
                8'h6:   segments = 7'h7D;
                8'h7:   segments = 7'h07;
                8'h8:   segments = 7'h7F;
                8'h9:   segments = 7'h67;
                8'hA:   segments = 7'h77;
                8'hB:   segments = 7'h7C;
                8'hC:   segments = 7'h39;
                8'hD:   segments = 7'h5E;
                8'hE:   segments = 7'h79;
                8'hF:   segments = 7'h71;
                default: segments = 7'h7f;
            endcase
       end

    assign out = ~segments;
endmodule


module hexdisplay(input [31:0] in, output [41:0] hexleds);
    hexLEDDriver segment0(.value((in & 32'h0000_000F)),       .out(hexleds[6:0]));
    hexLEDDriver segment1(.value((in & 32'h0000_00F0) >> 4),  .out(hexleds[13:7]));
    hexLEDDriver segment2(.value((in & 32'h0000_0F00) >> 8),  .out(hexleds[20:14]));
    hexLEDDriver segment3(.value((in & 32'h0000_F000) >> 12), .out(hexleds[27:21]));
    hexLEDDriver segment4(.value((in & 32'h000F_0000) >> 16), .out(hexleds[34:28]));
    hexLEDDriver segment5(.value((in & 32'h00F0_0000) >> 20), .out(hexleds[41:35]));
endmodule

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module Top(

	//////////// CLOCK //////////
	input					CLOCK_50,
	//input					CLOCK2_50,
	//input					CLOCK3_50,
	//input					CLOCK4_50,

	//////////// SEG7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,

	//////////// KEY //////////
	input		     [3:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR

	//////////// SW //////////
	//input		     [9:0]		SW,

	//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	//inout		    [35:0]		GPIO_0,

	//////////// GPIO_1, GPIO_1 connect to GPIO Default //////////
	//inout		    [35:0]		GPIO_1
);


//=======================================================
//  REG/WIRE declarations
//=======================================================

reg [63:0] counter;
wire CLOCK_5;
wire reset;
wire pll_locked;

reg [6:0]  hex0;
reg [6:0]  hex1;
reg [6:0]  hex2;
reg [6:0]  hex3;
reg [6:0]  hex4;
reg [6:0]  hex5;
reg [31:0] hexleds;


//=======================================================
//  Structural coding
//=======================================================

pll10MHz pll_10(.refclk(CLOCK_50), .rst(reset), .outclk_0(CLOCK_5), .locked(pll_locked));
assign reset  = 0;
assign LEDR[9] = pll_locked;


always @(posedge CLOCK_5)
    begin
        counter <= counter + 1;
        hexleds <= counter[51:20];
    end


//hexdisplay display(.x(32'h123456), .hexleds({HEX5, HEX4, HEX3, HEX2, HEX1, HEX0}));
hexdisplay display(.in(hexleds), .hexleds({HEX5, HEX4, HEX3, HEX2, HEX1, HEX0}));

assign LEDR[0]  = ~KEY[0];
assign LEDR[1]  = ~KEY[1];
assign LEDR[2]  = ~KEY[2];
assign LEDR[3]  = ~KEY[3];

//assign GPIO_0 = 0;
//assign GPIO_1 = 0;

endmodule
